module ui

interface DrawDevice {
}
