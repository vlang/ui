module editor
