module main

import ui

const (
	win_width = 250
	win_height = 250
)

struct App {
mut:
	hor_slider  &ui.Slider
	vert_slider &ui.Slider
	window      &ui.Window
}

fn main() {
	mut app := &App{}
	window := ui.window({
		width: win_width
		height: win_height
		title: 'Slider Example'
		user_ptr: app
	}, [
		ui.row({
			stretch: true
			alignment: .center
			margin: ui.MarginConfig{5,5,5,5}
			spacing: 10
		}, [
			ui.slider({
				width: 20
				height: 200
				orientation: .vertical
				max: 100
				val: 0
				on_value_changed: on_vert_value_changed
			}) as ui.IWidgeter,
			ui.slider({
				width: 200
				height: 20
				orientation: .horizontal
				max: 100
				val: 0
				on_value_changed: on_hor_value_changed
			})
		]) as ui.IWidgeter
	])
	app.window = window
	ui.run(window)
}

fn on_hor_value_changed(app mut App) {
	//app.vert_slider.val = app.hor_slider.val
}

fn on_vert_value_changed(app mut App) {
	//app.hor_slider.val = app.vert_slider.val
}
