module component

import ui
import gx

type ColorButtonFn = fn (b &ColorButtonComponent)

struct ColorButtonComponent {
pub mut:
	widget     &ui.Button
	bg_color   gx.Color = gx.white
	ctrl_mode  bool
	on_click   ColorButtonFn
	on_changed ColorButtonFn
}

[params]
pub struct ColorButtonParams {
	id           string
	text         string
	height       int
	width        int
	z_index      int
	tooltip      string
	tooltip_side ui.Side = .top
	radius       f64     = .25
	padding      f64
	bg_color     &gx.Color = 0
	ctrl_mode    bool
	on_click     ColorButtonFn
	on_changed   ColorButtonFn
}

pub fn colorbutton(c ColorButtonParams) &ui.Button {
	mut b := &ui.Button{
		id: c.id
		width_: c.width
		height_: c.height
		z_index: c.z_index
		bg_color: c.bg_color
		theme_cfg: ui.no_theme
		tooltip: ui.TooltipMessage{c.tooltip, c.tooltip_side}
		onclick: colorbutton_click
		radius: f32(c.radius)
		padding: f32(c.padding)
		ui: 0
	}
	cbc := &ColorButtonComponent{
		widget: b
		ctrl_mode: c.ctrl_mode
		on_click: c.on_click
		on_changed: c.on_changed
	}
	if b.bg_color == 0 {
		b.bg_color = &cbc.bg_color
	}
	ui.component_connect(cbc, b)
	return b
}

// component access
pub fn colorbutton_component(w ui.ComponentChild) &ColorButtonComponent {
	return &ColorButtonComponent(w.component)
}

pub fn colorbutton_component_from_id(w ui.Window, id string) &ColorButtonComponent {
	return colorbutton_component(w.button(id))
}

fn colorbutton_click(a voidptr, mut b ui.Button) {
	cbc := colorbutton_component(b)
	// println("here $cbc.ctrl_mode $b.ui.keymods")
	if !cbc.ctrl_mode || ui.ctrl_key(b.ui.keymods) {
		colorbox_subwindow_connect(b.ui.window, b.bg_color, cbc, true)
		// move only if s.x and s.y == 0 first use
		mut s := b.ui.window.subwindow(colorbox_subwindow_id)
		if s.x == 0 && s.y == 0 {
			w, h := b.size()
			s.set_pos(b.x + w / 2, b.y + h / 2)
			s.update_layout()
		}
	} else if cbc.ctrl_mode {
		mut s := b.ui.window.subwindow(colorbox_subwindow_id)
		if s.is_visible() {
			colorbox_subwindow_connect(b.ui.window, b.bg_color, cbc, false)
		}
	}
	// on_click initialization if necessary
	if cbc.on_click != ColorButtonFn(0) {
		cbc.on_click(cbc)
	}
}
