module ui

import gx

pub enum Cursor {
	hand
	arrow
	ibeam
}

pub fn draw_text(x, y int, s string, cfg gx.TextCfg) {

}

pub fn draw_text_def(x, y int, s string) {
}
