// Copyright (c) 2020-2022 Alexander Medvednikov. All rights reserved.
// Use of this source code is governed by a GPL license
// that can be found in the LICENSE file.
module ui

// This provides user defined shortcut actions (see grid and grid_data as a use case)
pub type ShortcutFn = fn (context voidptr)

pub type KeyShortcuts = map[int]Shortcut
pub type CharShortcuts = map[string]Shortcut

pub struct Shortcut {
pub mut:
	mods   KeyMod
	key_fn ShortcutFn
}

pub fn char_shortcut(e KeyEvent, shortcuts CharShortcuts, context voidptr) {
	// weirdly when .ctrl modifier the codepoint is differently interpreted
	s := if e.mods == .ctrl { rune(96 + e.codepoint).str() } else { utf32_to_str(e.codepoint) }
	if s in shortcuts {
		sc := shortcuts[s]
		if has_key_mods(e.mods, sc.mods) {
			sc.key_fn(context)
		}
	}
}

pub fn key_shortcut(e KeyEvent, shortcuts KeyShortcuts, context voidptr) {
	if int(e.key) in shortcuts {
		sc := shortcuts[int(e.key)]
		if has_key_mods(e.mods, sc.mods) {
			sc.key_fn(context)
		}
	}
}

pub interface Shortcutable {
	id string
mut:
	key_shortcuts KeyShortcuts
	char_shortcuts CharShortcuts
}

pub fn (mut s Shortcutable) add_char_shortcut(code string, mods KeyMod, key_fn ShortcutFn) {
	s.char_shortcuts[code] = Shortcut{
		mods: mods
		key_fn: key_fn
	}
}

pub fn (mut s Shortcutable) add_key_shortcut(code int, mods KeyMod, key_fn ShortcutFn) {
	s.key_shortcuts[code] = Shortcut{
		mods: mods
		key_fn: key_fn
	}
}

// BitMask

[flag]
pub enum KeyMod {
	shift //= 1 // (1<<0)
	ctrl //= 2 // (1<<1)
	alt //= 4 // (1<<2)
	super //= 8 // (1<<3)
}

pub enum KeyState {
	press = 1
	release = 0
	repeat = 2
}

pub struct KeyEvent {
pub:
	key       Key
	action    int
	code      int
	mods      KeyMod
	codepoint u32
}

// Copied from sapp/enums TODO alias?
pub enum Key {
	invalid = 0
	space = 32
	apostrophe = 39 // '
	comma = 44 // ,
	minus = 45 // -
	period = 46 // .
	slash = 47 // /
	_0 = 48
	_1 = 49
	_2 = 50
	_3 = 51
	_4 = 52
	_5 = 53
	_6 = 54
	_7 = 55
	_8 = 56
	_9 = 57
	semicolon = 59 // ;
	equal = 61 // =
	a = 65
	b = 66
	c = 67
	d = 68
	e = 69
	f = 70
	g = 71
	h = 72
	i = 73
	j = 74
	k = 75
	l = 76
	m = 77
	n = 78
	o = 79
	p = 80
	q = 81
	r = 82
	s = 83
	t = 84
	u = 85
	v = 86
	w = 87
	x = 88
	y = 89
	z = 90
	left_bracket = 91 // [
	backslash = 92 // \
	right_bracket = 93 // ]
	grave_accent = 96 // `
	world_1 = 161 // non-us #1
	world_2 = 162 // non-us #2
	escape = 256
	enter = 257
	tab = 258
	backspace = 259
	insert = 260
	delete = 261
	right = 262
	left = 263
	down = 264
	up = 265
	page_up = 266
	page_down = 267
	home = 268
	end = 269
	caps_lock = 280
	scroll_lock = 281
	num_lock = 282
	print_screen = 283
	pause = 284
	f1 = 290
	f2 = 291
	f3 = 292
	f4 = 293
	f5 = 294
	f6 = 295
	f7 = 296
	f8 = 297
	f9 = 298
	f10 = 299
	f11 = 300
	f12 = 301
	f13 = 302
	f14 = 303
	f15 = 304
	f16 = 305
	f17 = 306
	f18 = 307
	f19 = 308
	f20 = 309
	f21 = 310
	f22 = 311
	f23 = 312
	f24 = 313
	f25 = 314
	kp_0 = 320
	kp_1 = 321
	kp_2 = 322
	kp_3 = 323
	kp_4 = 324
	kp_5 = 325
	kp_6 = 326
	kp_7 = 327
	kp_8 = 328
	kp_9 = 329
	kp_decimal = 330
	kp_divide = 331
	kp_multiply = 332
	kp_subtract = 333
	kp_add = 334
	kp_enter = 335
	kp_equal = 336
	left_shift = 340
	left_control = 341
	left_alt = 342
	left_super = 343
	right_shift = 344
	right_control = 345
	right_alt = 346
	right_super = 347
	menu = 348
}

pub fn shift_key(mods KeyMod) bool {
	return int(mods) & 1 == 1
}

pub fn ctl_key(mods KeyMod) bool {
	return int(mods) & 2 == 2
}

pub fn alt_key(mods KeyMod) bool {
	return int(mods) & 4 == 4
}

pub fn super_key(mods KeyMod) bool {
	return int(mods) & 8 == 8
}

pub fn ctl_shift_key(mods KeyMod) bool {
	return int(mods) & 3 == 3
}

pub fn ctl_alt_key(mods KeyMod) bool {
	return int(mods) & 6 == 6
}

pub fn super_alt_key(mods KeyMod) bool {
	return int(mods) & 12 == 12
}

pub fn has_key_mods(mods KeyMod, opts KeyMod) bool {
	return int(mods) & int(opts) == int(opts)
}

// NB: to complete if useful
