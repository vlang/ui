module ui
const (
bytes_check_png_len = 3811
bytes_check_png = [ byte(
137), 80, 78, 71, 13, 10, 26, 10, 0, 0, 0, 13, 73, 72, 68, 82, 0, 0, 0, 16, 0, 0, 0, 16, 8, 6, 0, 0, 0, 31, 243, 255, 97, 0, 0, 0, 4, 103, 65, 77, 65, 0, 0, 177, 142, 124, 251, 81, 147, 0, 0, 0, 32, 99, 72, 82, 77, 0, 0, 135, 14, 0, 0, 140, 18, 0, 1, 10, 118, 0, 0, 124, 199, 0, 0, 108, 171, 0, 1, 10, 41, 0, 0, 60, 174, 0, 0, 22, 177, 136, 240, 182, 122, 0, 0, 10, 169, 105, 67, 67, 80, 73, 67, 67, 32, 80, 114, 111, 102, 105, 108, 101, 0, 0, 72, 199, 173, 150, 103, 84, 83, 217, 22, 199, 207, 189, 233, 141, 22, 64, 64, 74, 232, 189, 119, 144, 94, 67, 17, 164, 131, 168, 132, 36, 64, 40, 33, 36, 4, 20, 27, 34, 131, 35, 56, 22, 68, 68, 64, 29, 209, 65, 138, 130, 131, 82, 100, 16, 21, 11, 182, 65, 65, 193, 238, 128, 136, 128, 50, 78, 44, 216, 80, 51, 23, 120, 196, 153, 15, 239, 195, 91, 235, 237, 181, 118, 206, 111, 237, 181, 207, 62, 123, 223, 156, 179, 214, 31, 0, 242, 29, 6, 143, 151, 14, 203, 0, 144, 193, 205, 230, 135, 249, 121, 210, 98, 98, 227, 104, 184, 103, 0, 2, 48, 80, 0, 246, 64, 137, 193, 20, 240, 60, 66, 67, 131, 0, 98, 11, 235, 191, 237, 253, 16, 146, 141, 216, 109, 211, 217, 90, 224, 127, 51, 89, 22, 91, 192, 4, 0, 10, 69, 56, 145, 37, 96, 102, 32, 124, 10, 241, 46, 38, 143, 159, 13, 0, 138, 135, 196, 181, 115, 179, 121, 179, 92, 134, 176, 60, 31, 105, 16, 225, 186, 89, 78, 158, 231, 174, 89, 78, 156, 231, 91, 115, 57, 17, 97, 94, 8, 63, 3, 0, 79, 102, 48, 248, 201, 0, 144, 68, 72, 156, 150, 195, 76, 70, 234, 144, 145, 105, 129, 5, 151, 197, 225, 34, 236, 142, 176, 43, 51, 133, 193, 66, 56, 31, 97, 147, 140, 140, 204, 89, 62, 134, 176, 65, 226, 63, 234, 36, 255, 171, 102, 162, 164, 38, 131, 145, 44, 225, 249, 89, 230, 12, 239, 205, 17, 240, 210, 25, 107, 192, 255, 219, 50, 210, 133, 11, 103, 104, 35, 78, 78, 225, 251, 135, 205, 158, 55, 251, 221, 210, 50, 3, 37, 204, 77, 92, 26, 178, 192, 28, 214, 124, 79, 179, 156, 34, 244, 143, 92, 96, 166, 192, 43, 110, 129, 89, 12, 239, 64, 201, 222, 244, 165, 65, 11, 156, 196, 241, 165, 75, 234, 100, 211, 35, 22, 152, 159, 25, 38, 169, 207, 22, 248, 132, 47, 48, 131, 255, 253, 44, 97, 90, 164, 135, 228, 92, 54, 93, 82, 51, 47, 37, 34, 122, 129, 115, 56, 81, 75, 23, 88, 144, 22, 30, 248, 61, 199, 75, 18, 231, 11, 195, 36, 61, 39, 241, 125, 37, 51, 102, 8, 254, 49, 23, 135, 46, 201, 207, 78, 137, 240, 151, 204, 200, 248, 222, 27, 91, 16, 35, 233, 129, 197, 246, 246, 145, 196, 185, 145, 146, 28, 94, 182, 167, 164, 62, 47, 61, 84, 146, 207, 78, 247, 147, 196, 5, 57, 225, 146, 189, 217, 200, 101, 251, 190, 55, 84, 242, 125, 82, 25, 1, 161, 11, 12, 56, 32, 24, 48, 0, 51, 155, 189, 58, 123, 182, 97, 175, 76, 222, 26, 62, 39, 57, 37, 155, 230, 129, 188, 24, 54, 141, 206, 101, 154, 153, 208, 172, 44, 172, 44, 0, 152, 125, 127, 243, 127, 175, 232, 230, 220, 187, 130, 148, 101, 191, 199, 138, 144, 187, 230, 42, 18, 139, 197, 109, 223, 99, 254, 151, 0, 104, 113, 6, 128, 88, 249, 61, 166, 223, 0, 128, 212, 32, 0, 87, 30, 51, 133, 252, 156, 249, 24, 122, 246, 7, 3, 136, 64, 26, 200, 3, 101, 160, 142, 220, 31, 3, 96, 10, 172, 128, 29, 112, 6, 238, 192, 7, 4, 128, 16, 16, 1, 98, 193, 74, 192, 4, 41, 32, 3, 240, 65, 46, 88, 7, 54, 129, 34, 80, 2, 118, 130, 61, 160, 18, 28, 4, 135, 65, 29, 56, 14, 90, 64, 59, 232, 2, 231, 193, 101, 112, 29, 220, 2, 131, 224, 33, 24, 6, 99, 224, 37, 16, 129, 247, 96, 6, 130, 32, 28, 68, 129, 168, 144, 50, 164, 1, 233, 66, 198, 144, 21, 228, 0, 185, 66, 62, 80, 16, 20, 6, 197, 66, 9, 80, 50, 196, 133, 132, 208, 58, 104, 51, 84, 2, 149, 66, 149, 208, 33, 168, 30, 250, 21, 58, 13, 157, 135, 174, 66, 253, 208, 125, 104, 4, 154, 132, 222, 64, 159, 97, 20, 76, 134, 229, 97, 53, 88, 15, 54, 135, 29, 96, 15, 56, 16, 142, 128, 87, 192, 201, 112, 22, 156, 7, 23, 194, 219, 225, 10, 184, 6, 62, 6, 183, 193, 231, 225, 235, 240, 32, 60, 12, 191, 132, 167, 81, 0, 69, 66, 41, 162, 52, 81, 166, 40, 7, 148, 23, 42, 4, 21, 135, 74, 66, 241, 81, 27, 80, 197, 168, 114, 84, 13, 170, 9, 213, 137, 234, 69, 221, 70, 13, 163, 166, 80, 159, 208, 88, 52, 21, 77, 67, 155, 162, 157, 209, 254, 232, 72, 52, 19, 157, 133, 222, 128, 222, 134, 174, 68, 215, 161, 219, 208, 23, 209, 183, 209, 35, 104, 17, 250, 27, 134, 130, 81, 197, 24, 99, 156, 48, 116, 76, 12, 38, 25, 147, 139, 41, 194, 148, 99, 106, 49, 173, 152, 75, 152, 65, 204, 24, 230, 61, 22, 139, 85, 196, 234, 99, 237, 177, 254, 216, 88, 108, 42, 118, 45, 118, 27, 118, 63, 182, 25, 123, 14, 219, 143, 29, 197, 78, 227, 112, 56, 101, 156, 49, 206, 5, 23, 130, 99, 224, 178, 113, 69, 184, 125, 184, 99, 184, 179, 184, 1, 220, 24, 238, 35, 158, 132, 215, 192, 91, 225, 125, 241, 113, 120, 46, 190, 0, 95, 142, 111, 192, 119, 227, 7, 240, 227, 248, 25, 130, 12, 65, 151, 224, 68, 8, 33, 176, 8, 107, 8, 59, 8, 71, 8, 157, 132, 155, 132, 49, 194, 12, 81, 150, 168, 79, 116, 33, 70, 16, 83, 137, 155, 136, 21, 196, 38, 226, 37, 226, 35, 226, 91, 18, 137, 164, 69, 114, 36, 45, 35, 113, 72, 249, 164, 10, 210, 9, 210, 21, 210, 8, 233, 19, 89, 142, 108, 68, 246, 34, 199, 147, 133, 228, 237, 228, 163, 228, 115, 228, 251, 228, 183, 20, 10, 69, 143, 226, 78, 137, 163, 100, 83, 182, 83, 234, 41, 23, 40, 79, 40, 31, 165, 168, 82, 102, 82, 116, 41, 150, 212, 70, 169, 42, 169, 54, 169, 1, 169, 87, 210, 4, 105, 93, 105, 15, 233, 149, 210, 121, 210, 229, 210, 39, 165, 111, 74, 79, 201, 16, 100, 244, 100, 188, 100, 24, 50, 27, 100, 170, 100, 78, 203, 220, 149, 153, 150, 165, 202, 90, 202, 134, 200, 102, 200, 110, 147, 109, 144, 189, 42, 59, 33, 135, 147, 211, 147, 243, 145, 99, 201, 21, 202, 29, 150, 187, 32, 55, 74, 69, 81, 181, 169, 94, 84, 38, 117, 51, 245, 8, 245, 18, 117, 76, 30, 43, 175, 47, 79, 151, 79, 149, 47, 145, 63, 46, 223, 39, 47, 82, 144, 83, 176, 81, 136, 82, 88, 173, 80, 165, 112, 70, 97, 88, 17, 165, 168, 167, 72, 87, 76, 87, 220, 161, 216, 162, 56, 164, 248, 121, 145, 218, 34, 143, 69, 236, 69, 91, 23, 53, 45, 26, 88, 244, 65, 105, 177, 146, 187, 18, 91, 169, 88, 169, 89, 105, 80, 233, 179, 50, 77, 217, 71, 57, 77, 121, 151, 114, 187, 242, 99, 21, 180, 138, 145, 202, 50, 149, 92, 149, 3, 42, 151, 84, 166, 22, 203, 47, 118, 94, 204, 92, 92, 188, 184, 101, 241, 3, 85, 88, 213, 72, 53, 76, 117, 173, 234, 97, 213, 27, 170, 211, 106, 234, 106, 126, 106, 60, 181, 125, 106, 23, 212, 166, 212, 21, 213, 221, 213, 83, 213, 203, 212, 187, 213, 39, 53, 168, 26, 174, 26, 28, 141, 50, 141, 179, 26, 47, 104, 10, 52, 15, 90, 58, 173, 130, 118, 145, 38, 210, 84, 213, 244, 215, 20, 106, 30, 210, 236, 211, 156, 209, 210, 215, 138, 212, 42, 208, 106, 214, 122, 172, 77, 212, 118, 208, 78, 210, 46, 211, 238, 209, 22, 233, 104, 232, 4, 235, 172, 211, 105, 212, 121, 160, 75, 208, 117, 208, 77, 209, 221, 171, 219, 171, 251, 65, 79, 95, 47, 90, 111, 139, 94, 187, 222, 132, 190, 146, 62, 93, 63, 79, 191, 81, 255, 145, 1, 197, 192, 205, 32, 203, 160, 198, 224, 142, 33, 214, 208, 193, 48, 205, 112, 191, 225, 45, 35, 216, 200, 214, 40, 197, 168, 202, 232, 166, 49, 108, 108, 103, 204, 49, 222, 111, 220, 111, 130, 49, 113, 52, 225, 154, 212, 152, 220, 53, 37, 155, 122, 152, 230, 152, 54, 154, 142, 152, 41, 154, 5, 153, 21, 152, 181, 155, 189, 50, 215, 49, 143, 51, 223, 101, 222, 107, 254, 205, 194, 214, 34, 221, 226, 136, 197, 67, 75, 57, 203, 0, 203, 2, 203, 78, 203, 55, 86, 70, 86, 76, 171, 42, 171, 59, 214, 20, 107, 95, 235, 141, 214, 29, 214, 175, 109, 140, 109, 216, 54, 7, 108, 238, 217, 82, 109, 131, 109, 183, 216, 246, 216, 126, 181, 179, 183, 227, 219, 53, 217, 77, 218, 235, 216, 39, 216, 87, 219, 223, 117, 144, 119, 8, 117, 216, 230, 112, 197, 17, 227, 232, 233, 184, 209, 177, 203, 241, 147, 147, 157, 83, 182, 83, 139, 211, 95, 206, 166, 206, 105, 206, 13, 206, 19, 75, 244, 151, 176, 151, 28, 89, 50, 234, 162, 229, 194, 112, 57, 228, 50, 236, 74, 115, 77, 112, 253, 217, 117, 216, 77, 211, 141, 225, 86, 227, 246, 212, 93, 219, 157, 229, 94, 235, 62, 238, 97, 232, 145, 234, 113, 204, 227, 149, 167, 133, 39, 223, 179, 213, 243, 131, 151, 147, 215, 122, 175, 115, 222, 40, 111, 63, 239, 98, 239, 62, 31, 57, 159, 72, 159, 74, 159, 39, 190, 90, 190, 201, 190, 141, 190, 34, 63, 91, 191, 181, 126, 231, 252, 49, 254, 129, 254, 187, 252, 239, 210, 213, 232, 76, 122, 61, 93, 20, 96, 31, 176, 62, 224, 98, 32, 57, 48, 60, 176, 50, 240, 105, 144, 81, 16, 63, 168, 51, 24, 14, 14, 8, 222, 29, 252, 104, 169, 238, 82, 238, 210, 246, 16, 16, 66, 15, 217, 29, 242, 56, 84, 63, 52, 43, 244, 183, 101, 216, 101, 161, 203, 170, 150, 61, 15, 179, 12, 91, 23, 214, 27, 78, 13, 95, 21, 222, 16, 254, 62, 194, 51, 98, 71, 196, 195, 72, 131, 72, 97, 100, 79, 148, 116, 84, 124, 84, 125, 212, 135, 104, 239, 232, 210, 232, 225, 24, 243, 152, 245, 49, 215, 99, 85, 98, 57, 177, 29, 113, 184, 184, 168, 184, 218, 184, 233, 229, 62, 203, 247, 44, 31, 139, 183, 141, 47, 138, 31, 90, 161, 191, 98, 245, 138, 171, 43, 85, 86, 166, 175, 60, 179, 74, 122, 21, 99, 213, 201, 4, 76, 66, 116, 66, 67, 194, 23, 70, 8, 163, 134, 49, 157, 72, 79, 172, 78, 20, 49, 189, 152, 123, 153, 47, 89, 238, 172, 50, 214, 36, 219, 133, 93, 202, 30, 79, 114, 73, 42, 77, 154, 72, 118, 73, 222, 157, 60, 153, 226, 150, 82, 158, 50, 197, 241, 226, 84, 114, 94, 167, 250, 167, 30, 76, 253, 144, 22, 146, 118, 52, 77, 156, 30, 157, 222, 156, 129, 207, 72, 200, 56, 205, 149, 227, 166, 113, 47, 102, 170, 103, 174, 206, 236, 231, 25, 243, 138, 120, 195, 89, 78, 89, 123, 178, 68, 252, 64, 126, 173, 0, 18, 172, 16, 116, 100, 203, 35, 66, 231, 134, 208, 64, 248, 131, 112, 36, 199, 53, 167, 42, 231, 99, 110, 84, 238, 201, 213, 178, 171, 185, 171, 111, 172, 49, 90, 179, 117, 205, 120, 158, 111, 222, 47, 107, 209, 107, 153, 107, 123, 214, 105, 174, 219, 180, 110, 100, 189, 199, 250, 67, 27, 160, 13, 137, 27, 122, 54, 106, 111, 44, 220, 56, 150, 239, 151, 95, 183, 137, 184, 41, 109, 211, 239, 5, 22, 5, 165, 5, 239, 54, 71, 111, 238, 44, 84, 43, 204, 47, 28, 253, 193, 239, 135, 198, 34, 169, 34, 126, 209, 221, 45, 206, 91, 14, 254, 136, 254, 145, 243, 99, 223, 86, 235, 173, 251, 182, 126, 43, 102, 21, 95, 43, 177, 40, 41, 47, 249, 178, 141, 185, 237, 218, 79, 150, 63, 85, 252, 36, 222, 158, 180, 189, 111, 135, 221, 142, 3, 59, 177, 59, 185, 59, 135, 118, 185, 237, 170, 43, 149, 45, 205, 43, 29, 221, 29, 188, 187, 173, 140, 86, 86, 92, 246, 110, 207, 170, 61, 87, 203, 109, 202, 15, 238, 37, 238, 21, 238, 29, 174, 8, 170, 232, 216, 167, 179, 111, 231, 190, 47, 149, 41, 149, 131, 85, 158, 85, 205, 213, 170, 213, 91, 171, 63, 236, 103, 237, 31, 56, 224, 126, 160, 233, 160, 218, 193, 146, 131, 159, 127, 230, 252, 124, 239, 144, 223, 161, 182, 26, 189, 154, 242, 195, 216, 195, 57, 135, 159, 31, 137, 58, 210, 251, 139, 195, 47, 245, 181, 42, 181, 37, 181, 95, 143, 114, 143, 14, 215, 133, 213, 93, 172, 183, 175, 175, 111, 80, 109, 216, 209, 8, 55, 10, 27, 39, 143, 197, 31, 187, 117, 220, 251, 120, 71, 147, 105, 211, 161, 102, 197, 230, 146, 19, 224, 132, 240, 196, 139, 95, 19, 126, 29, 106, 9, 108, 233, 57, 233, 112, 178, 233, 148, 238, 169, 234, 86, 106, 107, 113, 27, 212, 182, 166, 77, 212, 158, 210, 62, 220, 17, 219, 209, 127, 58, 224, 116, 79, 167, 115, 103, 235, 111, 102, 191, 29, 237, 210, 236, 170, 58, 163, 112, 102, 71, 55, 177, 187, 176, 91, 124, 54, 239, 236, 244, 57, 222, 185, 169, 243, 201, 231, 71, 123, 86, 245, 60, 188, 16, 115, 225, 206, 197, 101, 23, 251, 46, 5, 94, 186, 114, 217, 247, 242, 133, 94, 143, 222, 179, 87, 92, 174, 116, 93, 117, 186, 122, 250, 154, 195, 181, 246, 235, 118, 215, 219, 110, 216, 222, 104, 253, 221, 246, 247, 214, 62, 187, 190, 182, 155, 246, 55, 59, 110, 57, 222, 234, 236, 95, 210, 223, 61, 224, 54, 112, 254, 182, 247, 237, 203, 119, 232, 119, 174, 15, 46, 29, 236, 31, 138, 28, 186, 119, 55, 254, 238, 240, 61, 214, 189, 137, 251, 233, 247, 95, 63, 200, 121, 48, 243, 48, 255, 17, 230, 81, 241, 99, 153, 199, 229, 79, 84, 159, 212, 252, 97, 248, 71, 243, 176, 221, 240, 153, 17, 239, 145, 27, 79, 195, 159, 62, 28, 101, 142, 190, 124, 38, 120, 246, 101, 172, 240, 57, 229, 121, 249, 184, 198, 120, 253, 132, 213, 68, 215, 164, 239, 228, 173, 23, 203, 95, 140, 189, 228, 189, 156, 153, 42, 250, 83, 246, 207, 234, 87, 6, 175, 78, 253, 229, 254, 215, 13, 81, 140, 104, 236, 53, 255, 181, 248, 205, 182, 183, 202, 111, 143, 190, 179, 121, 215, 51, 29, 58, 253, 228, 125, 198, 251, 153, 15, 197, 31, 149, 63, 214, 125, 114, 248, 212, 251, 57, 250, 243, 248, 76, 238, 23, 220, 151, 138, 175, 134, 95, 59, 191, 5, 126, 123, 36, 206, 16, 139, 121, 12, 62, 99, 78, 10, 160, 16, 135, 147, 146, 0, 120, 115, 20, 0, 74, 44, 0, 84, 68, 55, 19, 151, 207, 235, 227, 57, 131, 230, 53, 253, 28, 129, 255, 198, 243, 26, 122, 206, 236, 0, 104, 66, 150, 89, 41, 52, 43, 249, 78, 34, 90, 90, 15, 209, 214, 148, 115, 0, 132, 32, 107, 132, 59, 128, 173, 173, 37, 254, 31, 19, 36, 89, 91, 205, 215, 146, 106, 4, 0, 167, 41, 22, 191, 201, 4, 128, 128, 248, 23, 63, 177, 120, 38, 84, 44, 254, 90, 141, 52, 123, 7, 128, 238, 137, 121, 93, 62, 107, 88, 68, 191, 55, 81, 207, 11, 106, 227, 6, 190, 229, 231, 255, 91, 29, 3, 240, 55, 74, 247, 10, 138, 238, 200, 114, 131, 0, 0, 0, 9, 112, 72, 89, 115, 0, 0, 14, 196, 0, 0, 14, 196, 1, 149, 43, 14, 27, 0, 0, 2, 4, 105, 84, 88, 116, 88, 77, 76, 58, 99, 111, 109, 46, 97, 100, 111, 98, 101, 46, 120, 109, 112, 0, 0, 0, 0, 0, 60, 120, 58, 120, 109, 112, 109, 101, 116, 97, 32, 120, 109, 108, 110, 115, 58, 120, 61, 34, 97, 100, 111, 98, 101, 58, 110, 115, 58, 109, 101, 116, 97, 47, 34, 32, 120, 58, 120, 109, 112, 116, 107, 61, 34, 88, 77, 80, 32, 67, 111, 114, 101, 32, 53, 46, 52, 46, 48, 34, 62, 10, 32, 32, 32, 60, 114, 100, 102, 58, 82, 68, 70, 32, 120, 109, 108, 110, 115, 58, 114, 100, 102, 61, 34, 104, 116, 116, 112, 58, 47, 47, 119, 119, 119, 46, 119, 51, 46, 111, 114, 103, 47, 49, 57, 57, 57, 47, 48, 50, 47, 50, 50, 45, 114, 100, 102, 45, 115, 121, 110, 116, 97, 120, 45, 110, 115, 35, 34, 62, 10, 32, 32, 32, 32, 32, 32, 60, 114, 100, 102, 58, 68, 101, 115, 99, 114, 105, 112, 116, 105, 111, 110, 32, 114, 100, 102, 58, 97, 98, 111, 117, 116, 61, 34, 34, 10, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 120, 109, 108, 110, 115, 58, 101, 120, 105, 102, 61, 34, 104, 116, 116, 112, 58, 47, 47, 110, 115, 46, 97, 100, 111, 98, 101, 46, 99, 111, 109, 47, 101, 120, 105, 102, 47, 49, 46, 48, 47, 34, 10, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 120, 109, 108, 110, 115, 58, 116, 105, 102, 102, 61, 34, 104, 116, 116, 112, 58, 47, 47, 110, 115, 46, 97, 100, 111, 98, 101, 46, 99, 111, 109, 47, 116, 105, 102, 102, 47, 49, 46, 48, 47, 34, 62, 10, 32, 32, 32, 32, 32, 32, 32, 32, 32, 60, 101, 120, 105, 102, 58, 80, 105, 120, 101, 108, 89, 68, 105, 109, 101, 110, 115, 105, 111, 110, 62, 49, 53, 50, 60, 47, 101, 120, 105, 102, 58, 80, 105, 120, 101, 108, 89, 68, 105, 109, 101, 110, 115, 105, 111, 110, 62, 10, 32, 32, 32, 32, 32, 32, 32, 32, 32, 60, 101, 120, 105, 102, 58, 80, 105, 120, 101, 108, 88, 68, 105, 109, 101, 110, 115, 105, 111, 110, 62, 50, 50, 48, 60, 47, 101, 120, 105, 102, 58, 80, 105, 120, 101, 108, 88, 68, 105, 109, 101, 110, 115, 105, 111, 110, 62, 10, 32, 32, 32, 32, 32, 32, 32, 32, 32, 60, 116, 105, 102, 102, 58, 79, 114, 105, 101, 110, 116, 97, 116, 105, 111, 110, 62, 49, 60, 47, 116, 105, 102, 102, 58, 79, 114, 105, 101, 110, 116, 97, 116, 105, 111, 110, 62, 10, 32, 32, 32, 32, 32, 32, 60, 47, 114, 100, 102, 58, 68, 101, 115, 99, 114, 105, 112, 116, 105, 111, 110, 62, 10, 32, 32, 32, 60, 47, 114, 100, 102, 58, 82, 68, 70, 62, 10, 60, 47, 120, 58, 120, 109, 112, 109, 101, 116, 97, 62, 10, 233, 63, 32, 177, 0, 0, 1, 148, 73, 68, 65, 84, 56, 79, 149, 147, 177, 175, 193, 80, 24, 197, 207, 171, 65, 98, 40, 18, 36, 54, 131, 201, 102, 53, 8, 179, 197, 98, 105, 68, 24, 108, 93, 25, 76, 254, 2, 137, 69, 194, 210, 196, 42, 86, 210, 177, 145, 144, 24, 172, 6, 131, 8, 131, 16, 34, 97, 161, 232, 115, 63, 183, 120, 201, 243, 94, 253, 146, 38, 223, 57, 105, 79, 239, 185, 183, 253, 50, 110, 224, 3, 142, 199, 35, 42, 149, 10, 6, 131, 1, 36, 73, 194, 199, 1, 173, 86, 11, 181, 90, 141, 102, 81, 20, 33, 208, 100, 145, 217, 108, 134, 102, 179, 201, 21, 16, 141, 70, 173, 7, 92, 175, 87, 52, 26, 13, 28, 14, 7, 210, 126, 191, 31, 153, 76, 198, 122, 64, 183, 219, 69, 191, 223, 231, 10, 200, 231, 243, 240, 122, 189, 214, 2, 86, 171, 21, 20, 69, 225, 10, 136, 199, 227, 116, 49, 254, 13, 184, 92, 46, 180, 244, 205, 102, 67, 218, 227, 241, 208, 219, 77, 40, 96, 191, 223, 211, 141, 191, 209, 235, 245, 160, 105, 26, 87, 64, 54, 155, 165, 254, 38, 2, 59, 146, 84, 42, 133, 66, 161, 128, 237, 118, 203, 237, 59, 187, 221, 14, 245, 122, 29, 231, 243, 153, 116, 36, 18, 65, 34, 145, 160, 217, 196, 166, 235, 122, 249, 116, 58, 97, 185, 92, 98, 177, 88, 32, 22, 139, 65, 16, 238, 205, 88, 248, 104, 52, 162, 217, 237, 118, 163, 84, 42, 193, 229, 114, 145, 54, 17, 146, 201, 36, 31, 65, 187, 108, 110, 214, 112, 56, 68, 167, 211, 161, 153, 145, 78, 167, 17, 8, 4, 184, 122, 98, 107, 183, 219, 229, 233, 116, 138, 249, 124, 78, 198, 120, 60, 134, 211, 233, 164, 47, 110, 189, 94, 147, 23, 14, 135, 33, 203, 242, 99, 101, 175, 208, 167, 204, 186, 22, 139, 69, 76, 38, 19, 110, 63, 113, 56, 28, 168, 86, 171, 8, 6, 131, 220, 249, 9, 69, 178, 94, 172, 159, 207, 231, 35, 243, 21, 246, 195, 188, 123, 152, 241, 88, 19, 235, 199, 86, 97, 183, 219, 185, 3, 132, 66, 33, 58, 161, 63, 97, 21, 94, 81, 85, 213, 184, 109, 172, 145, 203, 229, 140, 91, 37, 238, 190, 195, 48, 190, 1, 231, 96, 208, 15, 105, 22, 68, 122, 0, 0, 0, 0, 73, 69, 78, 68, 174, 66, 96, 130, 
]!!)
