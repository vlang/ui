module ui

interface WidgetThemeStyle {
mut:
	id string
	theme_style string
}

pub fn (l Widget) update_them_style() {

}

pub fn (l Layout) update_them_style() {

}