module webview

// TODO: get dynamic username and latest/fixed version
// #flag windows -I C:\Users\USERNAME\.nuget\packages\microsoft.web.webview2\VERSION\build\native\include
#include <WebView2.h>

fn create_windows_web_view(url string, title string) {

}
