// v ui public consts
module ui

public const (
  font_dir = []string{
    r'c:\windows\fonts\arial.ttf',
    
  }
  
  // error massages
  img_notfound = 'Image file not found.'
  font_notfound = 'System font file not found.'
  glfw_notinstalled = 'glfw not installed.'
  freetype_notinstalled = 'freetype is not installed.'
  
  // default size
  default_font_size = 13
  default_height = 20
  
)
