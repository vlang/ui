module webview

#flag darwin -framework WebKit
#include "@VROOT/webview/webview_darwin.m"
